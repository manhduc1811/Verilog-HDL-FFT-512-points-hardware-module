module ROM_256(
	input clk,
	input in_valid,
	input rst_n,
	output reg [23:0] w_r,
	output reg [23:0] w_i,
	output reg[1:0] state
);
////////////////////////////////////////////
// Internal signals
reg       valid,next_valid;
reg [9:0] count,next_count;
////////////////////////////////////////////
// Next state logic
always @(*) begin
    if(in_valid || valid)next_count = count + 1;
    else next_count = count;
    
    if (count<10'd256) 
        state = 2'd0;
    else if (count >= 10'd256 && count < 10'd512)
        state = 2'd1;
    else if (count >= 10'd512 && count < 10'd768)
        state = 2'd2;
    else state = 2'd3;

	case(count)
	10'd512: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 000000000000000000000000;
	 next_valid = 1'b1;
	 end
	10'd513: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111101;
	 next_valid = 1'b1;
	 end
	10'd514: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111111010;
	 next_valid = 1'b1;
	 end
	10'd515: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110111;
	 next_valid = 1'b1;
	 end
	10'd516: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110011;
	 next_valid = 1'b1;
	 end
	10'd517: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 111111111111111111110000;
	 next_valid = 1'b1;
	 end
	10'd518: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101101;
	 next_valid = 1'b1;
	 end
	10'd519: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111101010;
	 next_valid = 1'b1;
	 end
	10'd520: begin 
	 w_r = 24'b 000000000000000011111111;
	 w_i = 24'b 111111111111111111100111;
	 next_valid = 1'b1;
	 end
	10'd521: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111100100;
	 next_valid = 1'b1;
	 end
	10'd522: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111100001;
	 next_valid = 1'b1;
	 end
	10'd523: begin 
	 w_r = 24'b 000000000000000011111110;
	 w_i = 24'b 111111111111111111011110;
	 next_valid = 1'b1;
	 end
	10'd524: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111011010;
	 next_valid = 1'b1;
	 end
	10'd525: begin 
	 w_r = 24'b 000000000000000011111101;
	 w_i = 24'b 111111111111111111010111;
	 next_valid = 1'b1;
	 end
	10'd526: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010100;
	 next_valid = 1'b1;
	 end
	10'd527: begin 
	 w_r = 24'b 000000000000000011111100;
	 w_i = 24'b 111111111111111111010001;
	 next_valid = 1'b1;
	 end
	10'd528: begin 
	 w_r = 24'b 000000000000000011111011;
	 w_i = 24'b 111111111111111111001110;
	 next_valid = 1'b1;
	 end
	10'd529: begin 
	 w_r = 24'b 000000000000000011111010;
	 w_i = 24'b 111111111111111111001011;
	 next_valid = 1'b1;
	 end
	10'd530: begin 
	 w_r = 24'b 000000000000000011111010;
	 w_i = 24'b 111111111111111111001000;
	 next_valid = 1'b1;
	 end
	10'd531: begin 
	 w_r = 24'b 000000000000000011111001;
	 w_i = 24'b 111111111111111111000101;
	 next_valid = 1'b1;
	 end
	10'd532: begin 
	 w_r = 24'b 000000000000000011111000;
	 w_i = 24'b 111111111111111111000010;
	 next_valid = 1'b1;
	 end
	10'd533: begin 
	 w_r = 24'b 000000000000000011111000;
	 w_i = 24'b 111111111111111110111111;
	 next_valid = 1'b1;
	 end
	10'd534: begin 
	 w_r = 24'b 000000000000000011110111;
	 w_i = 24'b 111111111111111110111100;
	 next_valid = 1'b1;
	 end
	10'd535: begin 
	 w_r = 24'b 000000000000000011110110;
	 w_i = 24'b 111111111111111110111001;
	 next_valid = 1'b1;
	 end
	10'd536: begin 
	 w_r = 24'b 000000000000000011110101;
	 w_i = 24'b 111111111111111110110110;
	 next_valid = 1'b1;
	 end
	10'd537: begin 
	 w_r = 24'b 000000000000000011110100;
	 w_i = 24'b 111111111111111110110011;
	 next_valid = 1'b1;
	 end
	10'd538: begin 
	 w_r = 24'b 000000000000000011110011;
	 w_i = 24'b 111111111111111110110000;
	 next_valid = 1'b1;
	 end
	10'd539: begin 
	 w_r = 24'b 000000000000000011110010;
	 w_i = 24'b 111111111111111110101101;
	 next_valid = 1'b1;
	 end
	10'd540: begin 
	 w_r = 24'b 000000000000000011110001;
	 w_i = 24'b 111111111111111110101010;
	 next_valid = 1'b1;
	 end
	10'd541: begin 
	 w_r = 24'b 000000000000000011110000;
	 w_i = 24'b 111111111111111110100111;
	 next_valid = 1'b1;
	 end
	10'd542: begin 
	 w_r = 24'b 000000000000000011101111;
	 w_i = 24'b 111111111111111110100100;
	 next_valid = 1'b1;
	 end
	10'd543: begin 
	 w_r = 24'b 000000000000000011101110;
	 w_i = 24'b 111111111111111110100001;
	 next_valid = 1'b1;
	 end
	10'd544: begin 
	 w_r = 24'b 000000000000000011101101;
	 w_i = 24'b 111111111111111110011110;
	 next_valid = 1'b1;
	 end
	10'd545: begin 
	 w_r = 24'b 000000000000000011101011;
	 w_i = 24'b 111111111111111110011011;
	 next_valid = 1'b1;
	 end
	10'd546: begin 
	 w_r = 24'b 000000000000000011101010;
	 w_i = 24'b 111111111111111110011000;
	 next_valid = 1'b1;
	 end
	10'd547: begin 
	 w_r = 24'b 000000000000000011101001;
	 w_i = 24'b 111111111111111110010101;
	 next_valid = 1'b1;
	 end
	10'd548: begin 
	 w_r = 24'b 000000000000000011100111;
	 w_i = 24'b 111111111111111110010011;
	 next_valid = 1'b1;
	 end
	10'd549: begin 
	 w_r = 24'b 000000000000000011100110;
	 w_i = 24'b 111111111111111110010000;
	 next_valid = 1'b1;
	 end
	10'd550: begin 
	 w_r = 24'b 000000000000000011100101;
	 w_i = 24'b 111111111111111110001101;
	 next_valid = 1'b1;
	 end
	10'd551: begin 
	 w_r = 24'b 000000000000000011100011;
	 w_i = 24'b 111111111111111110001010;
	 next_valid = 1'b1;
	 end
	10'd552: begin 
	 w_r = 24'b 000000000000000011100010;
	 w_i = 24'b 111111111111111110000111;
	 next_valid = 1'b1;
	 end
	10'd553: begin 
	 w_r = 24'b 000000000000000011100000;
	 w_i = 24'b 111111111111111110000101;
	 next_valid = 1'b1;
	 end
	10'd554: begin 
	 w_r = 24'b 000000000000000011011111;
	 w_i = 24'b 111111111111111110000010;
	 next_valid = 1'b1;
	 end
	10'd555: begin 
	 w_r = 24'b 000000000000000011011101;
	 w_i = 24'b 111111111111111101111111;
	 next_valid = 1'b1;
	 end
	10'd556: begin 
	 w_r = 24'b 000000000000000011011100;
	 w_i = 24'b 111111111111111101111100;
	 next_valid = 1'b1;
	 end
	10'd557: begin 
	 w_r = 24'b 000000000000000011011010;
	 w_i = 24'b 111111111111111101111010;
	 next_valid = 1'b1;
	 end
	10'd558: begin 
	 w_r = 24'b 000000000000000011011000;
	 w_i = 24'b 111111111111111101110111;
	 next_valid = 1'b1;
	 end
	10'd559: begin 
	 w_r = 24'b 000000000000000011010111;
	 w_i = 24'b 111111111111111101110100;
	 next_valid = 1'b1;
	 end
	10'd560: begin 
	 w_r = 24'b 000000000000000011010101;
	 w_i = 24'b 111111111111111101110010;
	 next_valid = 1'b1;
	 end
	10'd561: begin 
	 w_r = 24'b 000000000000000011010011;
	 w_i = 24'b 111111111111111101101111;
	 next_valid = 1'b1;
	 end
	10'd562: begin 
	 w_r = 24'b 000000000000000011010001;
	 w_i = 24'b 111111111111111101101101;
	 next_valid = 1'b1;
	 end
	10'd563: begin 
	 w_r = 24'b 000000000000000011001111;
	 w_i = 24'b 111111111111111101101010;
	 next_valid = 1'b1;
	 end
	10'd564: begin 
	 w_r = 24'b 000000000000000011001110;
	 w_i = 24'b 111111111111111101101000;
	 next_valid = 1'b1;
	 end
	10'd565: begin 
	 w_r = 24'b 000000000000000011001100;
	 w_i = 24'b 111111111111111101100101;
	 next_valid = 1'b1;
	 end
	10'd566: begin 
	 w_r = 24'b 000000000000000011001010;
	 w_i = 24'b 111111111111111101100011;
	 next_valid = 1'b1;
	 end
	10'd567: begin 
	 w_r = 24'b 000000000000000011001000;
	 w_i = 24'b 111111111111111101100000;
	 next_valid = 1'b1;
	 end
	10'd568: begin 
	 w_r = 24'b 000000000000000011000110;
	 w_i = 24'b 111111111111111101011110;
	 next_valid = 1'b1;
	 end
	10'd569: begin 
	 w_r = 24'b 000000000000000011000100;
	 w_i = 24'b 111111111111111101011011;
	 next_valid = 1'b1;
	 end
	10'd570: begin 
	 w_r = 24'b 000000000000000011000010;
	 w_i = 24'b 111111111111111101011001;
	 next_valid = 1'b1;
	 end
	10'd571: begin 
	 w_r = 24'b 000000000000000011000000;
	 w_i = 24'b 111111111111111101010110;
	 next_valid = 1'b1;
	 end
	10'd572: begin 
	 w_r = 24'b 000000000000000010111110;
	 w_i = 24'b 111111111111111101010100;
	 next_valid = 1'b1;
	 end
	10'd573: begin 
	 w_r = 24'b 000000000000000010111100;
	 w_i = 24'b 111111111111111101010010;
	 next_valid = 1'b1;
	 end
	10'd574: begin 
	 w_r = 24'b 000000000000000010111001;
	 w_i = 24'b 111111111111111101001111;
	 next_valid = 1'b1;
	 end
	10'd575: begin 
	 w_r = 24'b 000000000000000010110111;
	 w_i = 24'b 111111111111111101001101;
	 next_valid = 1'b1;
	 end
	10'd576: begin 
	 w_r = 24'b 000000000000000010110101;
	 w_i = 24'b 111111111111111101001011;
	 next_valid = 1'b1;
	 end
	10'd577: begin 
	 w_r = 24'b 000000000000000010110011;
	 w_i = 24'b 111111111111111101001001;
	 next_valid = 1'b1;
	 end
	10'd578: begin 
	 w_r = 24'b 000000000000000010110001;
	 w_i = 24'b 111111111111111101000111;
	 next_valid = 1'b1;
	 end
	10'd579: begin 
	 w_r = 24'b 000000000000000010101110;
	 w_i = 24'b 111111111111111101000100;
	 next_valid = 1'b1;
	 end
	10'd580: begin 
	 w_r = 24'b 000000000000000010101100;
	 w_i = 24'b 111111111111111101000010;
	 next_valid = 1'b1;
	 end
	10'd581: begin 
	 w_r = 24'b 000000000000000010101010;
	 w_i = 24'b 111111111111111101000000;
	 next_valid = 1'b1;
	 end
	10'd582: begin 
	 w_r = 24'b 000000000000000010100111;
	 w_i = 24'b 111111111111111100111110;
	 next_valid = 1'b1;
	 end
	10'd583: begin 
	 w_r = 24'b 000000000000000010100101;
	 w_i = 24'b 111111111111111100111100;
	 next_valid = 1'b1;
	 end
	10'd584: begin 
	 w_r = 24'b 000000000000000010100010;
	 w_i = 24'b 111111111111111100111010;
	 next_valid = 1'b1;
	 end
	10'd585: begin 
	 w_r = 24'b 000000000000000010100000;
	 w_i = 24'b 111111111111111100111000;
	 next_valid = 1'b1;
	 end
	10'd586: begin 
	 w_r = 24'b 000000000000000010011101;
	 w_i = 24'b 111111111111111100110110;
	 next_valid = 1'b1;
	 end
	10'd587: begin 
	 w_r = 24'b 000000000000000010011011;
	 w_i = 24'b 111111111111111100110100;
	 next_valid = 1'b1;
	 end
	10'd588: begin 
	 w_r = 24'b 000000000000000010011000;
	 w_i = 24'b 111111111111111100110010;
	 next_valid = 1'b1;
	 end
	10'd589: begin 
	 w_r = 24'b 000000000000000010010110;
	 w_i = 24'b 111111111111111100110001;
	 next_valid = 1'b1;
	 end
	10'd590: begin 
	 w_r = 24'b 000000000000000010010011;
	 w_i = 24'b 111111111111111100101111;
	 next_valid = 1'b1;
	 end
	10'd591: begin 
	 w_r = 24'b 000000000000000010010001;
	 w_i = 24'b 111111111111111100101101;
	 next_valid = 1'b1;
	 end
	10'd592: begin 
	 w_r = 24'b 000000000000000010001110;
	 w_i = 24'b 111111111111111100101011;
	 next_valid = 1'b1;
	 end
	10'd593: begin 
	 w_r = 24'b 000000000000000010001100;
	 w_i = 24'b 111111111111111100101001;
	 next_valid = 1'b1;
	 end
	10'd594: begin 
	 w_r = 24'b 000000000000000010001001;
	 w_i = 24'b 111111111111111100101000;
	 next_valid = 1'b1;
	 end
	10'd595: begin 
	 w_r = 24'b 000000000000000010000110;
	 w_i = 24'b 111111111111111100100110;
	 next_valid = 1'b1;
	 end
	10'd596: begin 
	 w_r = 24'b 000000000000000010000100;
	 w_i = 24'b 111111111111111100100100;
	 next_valid = 1'b1;
	 end
	10'd597: begin 
	 w_r = 24'b 000000000000000010000001;
	 w_i = 24'b 111111111111111100100011;
	 next_valid = 1'b1;
	 end
	10'd598: begin 
	 w_r = 24'b 000000000000000001111110;
	 w_i = 24'b 111111111111111100100001;
	 next_valid = 1'b1;
	 end
	10'd599: begin 
	 w_r = 24'b 000000000000000001111011;
	 w_i = 24'b 111111111111111100100000;
	 next_valid = 1'b1;
	 end
	10'd600: begin 
	 w_r = 24'b 000000000000000001111001;
	 w_i = 24'b 111111111111111100011110;
	 next_valid = 1'b1;
	 end
	10'd601: begin 
	 w_r = 24'b 000000000000000001110110;
	 w_i = 24'b 111111111111111100011101;
	 next_valid = 1'b1;
	 end
	10'd602: begin 
	 w_r = 24'b 000000000000000001110011;
	 w_i = 24'b 111111111111111100011011;
	 next_valid = 1'b1;
	 end
	10'd603: begin 
	 w_r = 24'b 000000000000000001110000;
	 w_i = 24'b 111111111111111100011010;
	 next_valid = 1'b1;
	 end
	10'd604: begin 
	 w_r = 24'b 000000000000000001101101;
	 w_i = 24'b 111111111111111100011001;
	 next_valid = 1'b1;
	 end
	10'd605: begin 
	 w_r = 24'b 000000000000000001101011;
	 w_i = 24'b 111111111111111100010111;
	 next_valid = 1'b1;
	 end
	10'd606: begin 
	 w_r = 24'b 000000000000000001101000;
	 w_i = 24'b 111111111111111100010110;
	 next_valid = 1'b1;
	 end
	10'd607: begin 
	 w_r = 24'b 000000000000000001100101;
	 w_i = 24'b 111111111111111100010101;
	 next_valid = 1'b1;
	 end
	10'd608: begin 
	 w_r = 24'b 000000000000000001100010;
	 w_i = 24'b 111111111111111100010011;
	 next_valid = 1'b1;
	 end
	10'd609: begin 
	 w_r = 24'b 000000000000000001011111;
	 w_i = 24'b 111111111111111100010010;
	 next_valid = 1'b1;
	 end
	10'd610: begin 
	 w_r = 24'b 000000000000000001011100;
	 w_i = 24'b 111111111111111100010001;
	 next_valid = 1'b1;
	 end
	10'd611: begin 
	 w_r = 24'b 000000000000000001011001;
	 w_i = 24'b 111111111111111100010000;
	 next_valid = 1'b1;
	 end
	10'd612: begin 
	 w_r = 24'b 000000000000000001010110;
	 w_i = 24'b 111111111111111100001111;
	 next_valid = 1'b1;
	 end
	10'd613: begin 
	 w_r = 24'b 000000000000000001010011;
	 w_i = 24'b 111111111111111100001110;
	 next_valid = 1'b1;
	 end
	10'd614: begin 
	 w_r = 24'b 000000000000000001010000;
	 w_i = 24'b 111111111111111100001101;
	 next_valid = 1'b1;
	 end
	10'd615: begin 
	 w_r = 24'b 000000000000000001001101;
	 w_i = 24'b 111111111111111100001100;
	 next_valid = 1'b1;
	 end
	10'd616: begin 
	 w_r = 24'b 000000000000000001001010;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	10'd617: begin 
	 w_r = 24'b 000000000000000001000111;
	 w_i = 24'b 111111111111111100001010;
	 next_valid = 1'b1;
	 end
	10'd618: begin 
	 w_r = 24'b 000000000000000001000100;
	 w_i = 24'b 111111111111111100001001;
	 next_valid = 1'b1;
	 end
	10'd619: begin 
	 w_r = 24'b 000000000000000001000001;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	10'd620: begin 
	 w_r = 24'b 000000000000000000111110;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	10'd621: begin 
	 w_r = 24'b 000000000000000000111011;
	 w_i = 24'b 111111111111111100000111;
	 next_valid = 1'b1;
	 end
	10'd622: begin 
	 w_r = 24'b 000000000000000000111000;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	10'd623: begin 
	 w_r = 24'b 000000000000000000110101;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	10'd624: begin 
	 w_r = 24'b 000000000000000000110010;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	10'd625: begin 
	 w_r = 24'b 000000000000000000101111;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	10'd626: begin 
	 w_r = 24'b 000000000000000000101100;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	10'd627: begin 
	 w_r = 24'b 000000000000000000101001;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	10'd628: begin 
	 w_r = 24'b 000000000000000000100110;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	10'd629: begin 
	 w_r = 24'b 000000000000000000100010;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	10'd630: begin 
	 w_r = 24'b 000000000000000000011111;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	10'd631: begin 
	 w_r = 24'b 000000000000000000011100;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	10'd632: begin 
	 w_r = 24'b 000000000000000000011001;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	10'd633: begin 
	 w_r = 24'b 000000000000000000010110;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	10'd634: begin 
	 w_r = 24'b 000000000000000000010011;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	10'd635: begin 
	 w_r = 24'b 000000000000000000010000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd636: begin 
	 w_r = 24'b 000000000000000000001101;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd637: begin 
	 w_r = 24'b 000000000000000000001001;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd638: begin 
	 w_r = 24'b 000000000000000000000110;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd639: begin 
	 w_r = 24'b 000000000000000000000011;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd640: begin 
	 w_r = 24'b 000000000000000000000000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd641: begin 
	 w_r = 24'b 111111111111111111111101;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd642: begin 
	 w_r = 24'b 111111111111111111111010;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd643: begin 
	 w_r = 24'b 111111111111111111110111;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd644: begin 
	 w_r = 24'b 111111111111111111110011;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd645: begin 
	 w_r = 24'b 111111111111111111110000;
	 w_i = 24'b 111111111111111100000000;
	 next_valid = 1'b1;
	 end
	10'd646: begin 
	 w_r = 24'b 111111111111111111101101;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	10'd647: begin 
	 w_r = 24'b 111111111111111111101010;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	10'd648: begin 
	 w_r = 24'b 111111111111111111100111;
	 w_i = 24'b 111111111111111100000001;
	 next_valid = 1'b1;
	 end
	10'd649: begin 
	 w_r = 24'b 111111111111111111100100;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	10'd650: begin 
	 w_r = 24'b 111111111111111111100001;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	10'd651: begin 
	 w_r = 24'b 111111111111111111011110;
	 w_i = 24'b 111111111111111100000010;
	 next_valid = 1'b1;
	 end
	10'd652: begin 
	 w_r = 24'b 111111111111111111011010;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	10'd653: begin 
	 w_r = 24'b 111111111111111111010111;
	 w_i = 24'b 111111111111111100000011;
	 next_valid = 1'b1;
	 end
	10'd654: begin 
	 w_r = 24'b 111111111111111111010100;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	10'd655: begin 
	 w_r = 24'b 111111111111111111010001;
	 w_i = 24'b 111111111111111100000100;
	 next_valid = 1'b1;
	 end
	10'd656: begin 
	 w_r = 24'b 111111111111111111001110;
	 w_i = 24'b 111111111111111100000101;
	 next_valid = 1'b1;
	 end
	10'd657: begin 
	 w_r = 24'b 111111111111111111001011;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	10'd658: begin 
	 w_r = 24'b 111111111111111111001000;
	 w_i = 24'b 111111111111111100000110;
	 next_valid = 1'b1;
	 end
	10'd659: begin 
	 w_r = 24'b 111111111111111111000101;
	 w_i = 24'b 111111111111111100000111;
	 next_valid = 1'b1;
	 end
	10'd660: begin 
	 w_r = 24'b 111111111111111111000010;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	10'd661: begin 
	 w_r = 24'b 111111111111111110111111;
	 w_i = 24'b 111111111111111100001000;
	 next_valid = 1'b1;
	 end
	10'd662: begin 
	 w_r = 24'b 111111111111111110111100;
	 w_i = 24'b 111111111111111100001001;
	 next_valid = 1'b1;
	 end
	10'd663: begin 
	 w_r = 24'b 111111111111111110111001;
	 w_i = 24'b 111111111111111100001010;
	 next_valid = 1'b1;
	 end
	10'd664: begin 
	 w_r = 24'b 111111111111111110110110;
	 w_i = 24'b 111111111111111100001011;
	 next_valid = 1'b1;
	 end
	10'd665: begin 
	 w_r = 24'b 111111111111111110110011;
	 w_i = 24'b 111111111111111100001100;
	 next_valid = 1'b1;
	 end
	10'd666: begin 
	 w_r = 24'b 111111111111111110110000;
	 w_i = 24'b 111111111111111100001101;
	 next_valid = 1'b1;
	 end
	10'd667: begin 
	 w_r = 24'b 111111111111111110101101;
	 w_i = 24'b 111111111111111100001110;
	 next_valid = 1'b1;
	 end
	10'd668: begin 
	 w_r = 24'b 111111111111111110101010;
	 w_i = 24'b 111111111111111100001111;
	 next_valid = 1'b1;
	 end
	10'd669: begin 
	 w_r = 24'b 111111111111111110100111;
	 w_i = 24'b 111111111111111100010000;
	 next_valid = 1'b1;
	 end
	10'd670: begin 
	 w_r = 24'b 111111111111111110100100;
	 w_i = 24'b 111111111111111100010001;
	 next_valid = 1'b1;
	 end
	10'd671: begin 
	 w_r = 24'b 111111111111111110100001;
	 w_i = 24'b 111111111111111100010010;
	 next_valid = 1'b1;
	 end
	10'd672: begin 
	 w_r = 24'b 111111111111111110011110;
	 w_i = 24'b 111111111111111100010011;
	 next_valid = 1'b1;
	 end
	10'd673: begin 
	 w_r = 24'b 111111111111111110011011;
	 w_i = 24'b 111111111111111100010101;
	 next_valid = 1'b1;
	 end
	10'd674: begin 
	 w_r = 24'b 111111111111111110011000;
	 w_i = 24'b 111111111111111100010110;
	 next_valid = 1'b1;
	 end
	10'd675: begin 
	 w_r = 24'b 111111111111111110010101;
	 w_i = 24'b 111111111111111100010111;
	 next_valid = 1'b1;
	 end
	10'd676: begin 
	 w_r = 24'b 111111111111111110010011;
	 w_i = 24'b 111111111111111100011001;
	 next_valid = 1'b1;
	 end
	10'd677: begin 
	 w_r = 24'b 111111111111111110010000;
	 w_i = 24'b 111111111111111100011010;
	 next_valid = 1'b1;
	 end
	10'd678: begin 
	 w_r = 24'b 111111111111111110001101;
	 w_i = 24'b 111111111111111100011011;
	 next_valid = 1'b1;
	 end
	10'd679: begin 
	 w_r = 24'b 111111111111111110001010;
	 w_i = 24'b 111111111111111100011101;
	 next_valid = 1'b1;
	 end
	10'd680: begin 
	 w_r = 24'b 111111111111111110000111;
	 w_i = 24'b 111111111111111100011110;
	 next_valid = 1'b1;
	 end
	10'd681: begin 
	 w_r = 24'b 111111111111111110000101;
	 w_i = 24'b 111111111111111100100000;
	 next_valid = 1'b1;
	 end
	10'd682: begin 
	 w_r = 24'b 111111111111111110000010;
	 w_i = 24'b 111111111111111100100001;
	 next_valid = 1'b1;
	 end
	10'd683: begin 
	 w_r = 24'b 111111111111111101111111;
	 w_i = 24'b 111111111111111100100011;
	 next_valid = 1'b1;
	 end
	10'd684: begin 
	 w_r = 24'b 111111111111111101111100;
	 w_i = 24'b 111111111111111100100100;
	 next_valid = 1'b1;
	 end
	10'd685: begin 
	 w_r = 24'b 111111111111111101111010;
	 w_i = 24'b 111111111111111100100110;
	 next_valid = 1'b1;
	 end
	10'd686: begin 
	 w_r = 24'b 111111111111111101110111;
	 w_i = 24'b 111111111111111100101000;
	 next_valid = 1'b1;
	 end
	10'd687: begin 
	 w_r = 24'b 111111111111111101110100;
	 w_i = 24'b 111111111111111100101001;
	 next_valid = 1'b1;
	 end
	10'd688: begin 
	 w_r = 24'b 111111111111111101110010;
	 w_i = 24'b 111111111111111100101011;
	 next_valid = 1'b1;
	 end
	10'd689: begin 
	 w_r = 24'b 111111111111111101101111;
	 w_i = 24'b 111111111111111100101101;
	 next_valid = 1'b1;
	 end
	10'd690: begin 
	 w_r = 24'b 111111111111111101101101;
	 w_i = 24'b 111111111111111100101111;
	 next_valid = 1'b1;
	 end
	10'd691: begin 
	 w_r = 24'b 111111111111111101101010;
	 w_i = 24'b 111111111111111100110001;
	 next_valid = 1'b1;
	 end
	10'd692: begin 
	 w_r = 24'b 111111111111111101101000;
	 w_i = 24'b 111111111111111100110010;
	 next_valid = 1'b1;
	 end
	10'd693: begin 
	 w_r = 24'b 111111111111111101100101;
	 w_i = 24'b 111111111111111100110100;
	 next_valid = 1'b1;
	 end
	10'd694: begin 
	 w_r = 24'b 111111111111111101100011;
	 w_i = 24'b 111111111111111100110110;
	 next_valid = 1'b1;
	 end
	10'd695: begin 
	 w_r = 24'b 111111111111111101100000;
	 w_i = 24'b 111111111111111100111000;
	 next_valid = 1'b1;
	 end
	10'd696: begin 
	 w_r = 24'b 111111111111111101011110;
	 w_i = 24'b 111111111111111100111010;
	 next_valid = 1'b1;
	 end
	10'd697: begin 
	 w_r = 24'b 111111111111111101011011;
	 w_i = 24'b 111111111111111100111100;
	 next_valid = 1'b1;
	 end
	10'd698: begin 
	 w_r = 24'b 111111111111111101011001;
	 w_i = 24'b 111111111111111100111110;
	 next_valid = 1'b1;
	 end
	10'd699: begin 
	 w_r = 24'b 111111111111111101010110;
	 w_i = 24'b 111111111111111101000000;
	 next_valid = 1'b1;
	 end
	10'd700: begin 
	 w_r = 24'b 111111111111111101010100;
	 w_i = 24'b 111111111111111101000010;
	 next_valid = 1'b1;
	 end
	10'd701: begin 
	 w_r = 24'b 111111111111111101010010;
	 w_i = 24'b 111111111111111101000100;
	 next_valid = 1'b1;
	 end
	10'd702: begin 
	 w_r = 24'b 111111111111111101001111;
	 w_i = 24'b 111111111111111101000111;
	 next_valid = 1'b1;
	 end
	10'd703: begin 
	 w_r = 24'b 111111111111111101001101;
	 w_i = 24'b 111111111111111101001001;
	 next_valid = 1'b1;
	 end
	10'd704: begin 
	 w_r = 24'b 111111111111111101001011;
	 w_i = 24'b 111111111111111101001011;
	 next_valid = 1'b1;
	 end
	10'd705: begin 
	 w_r = 24'b 111111111111111101001001;
	 w_i = 24'b 111111111111111101001101;
	 next_valid = 1'b1;
	 end
	10'd706: begin 
	 w_r = 24'b 111111111111111101000111;
	 w_i = 24'b 111111111111111101001111;
	 next_valid = 1'b1;
	 end
	10'd707: begin 
	 w_r = 24'b 111111111111111101000100;
	 w_i = 24'b 111111111111111101010010;
	 next_valid = 1'b1;
	 end
	10'd708: begin 
	 w_r = 24'b 111111111111111101000010;
	 w_i = 24'b 111111111111111101010100;
	 next_valid = 1'b1;
	 end
	10'd709: begin 
	 w_r = 24'b 111111111111111101000000;
	 w_i = 24'b 111111111111111101010110;
	 next_valid = 1'b1;
	 end
	10'd710: begin 
	 w_r = 24'b 111111111111111100111110;
	 w_i = 24'b 111111111111111101011001;
	 next_valid = 1'b1;
	 end
	10'd711: begin 
	 w_r = 24'b 111111111111111100111100;
	 w_i = 24'b 111111111111111101011011;
	 next_valid = 1'b1;
	 end
	10'd712: begin 
	 w_r = 24'b 111111111111111100111010;
	 w_i = 24'b 111111111111111101011110;
	 next_valid = 1'b1;
	 end
	10'd713: begin 
	 w_r = 24'b 111111111111111100111000;
	 w_i = 24'b 111111111111111101100000;
	 next_valid = 1'b1;
	 end
	10'd714: begin 
	 w_r = 24'b 111111111111111100110110;
	 w_i = 24'b 111111111111111101100011;
	 next_valid = 1'b1;
	 end
	10'd715: begin 
	 w_r = 24'b 111111111111111100110100;
	 w_i = 24'b 111111111111111101100101;
	 next_valid = 1'b1;
	 end
	10'd716: begin 
	 w_r = 24'b 111111111111111100110010;
	 w_i = 24'b 111111111111111101101000;
	 next_valid = 1'b1;
	 end
	10'd717: begin 
	 w_r = 24'b 111111111111111100110001;
	 w_i = 24'b 111111111111111101101010;
	 next_valid = 1'b1;
	 end
	10'd718: begin 
	 w_r = 24'b 111111111111111100101111;
	 w_i = 24'b 111111111111111101101101;
	 next_valid = 1'b1;
	 end
	10'd719: begin 
	 w_r = 24'b 111111111111111100101101;
	 w_i = 24'b 111111111111111101101111;
	 next_valid = 1'b1;
	 end
	10'd720: begin 
	 w_r = 24'b 111111111111111100101011;
	 w_i = 24'b 111111111111111101110010;
	 next_valid = 1'b1;
	 end
	10'd721: begin 
	 w_r = 24'b 111111111111111100101001;
	 w_i = 24'b 111111111111111101110100;
	 next_valid = 1'b1;
	 end
	10'd722: begin 
	 w_r = 24'b 111111111111111100101000;
	 w_i = 24'b 111111111111111101110111;
	 next_valid = 1'b1;
	 end
	10'd723: begin 
	 w_r = 24'b 111111111111111100100110;
	 w_i = 24'b 111111111111111101111010;
	 next_valid = 1'b1;
	 end
	10'd724: begin 
	 w_r = 24'b 111111111111111100100100;
	 w_i = 24'b 111111111111111101111100;
	 next_valid = 1'b1;
	 end
	10'd725: begin 
	 w_r = 24'b 111111111111111100100011;
	 w_i = 24'b 111111111111111101111111;
	 next_valid = 1'b1;
	 end
	10'd726: begin 
	 w_r = 24'b 111111111111111100100001;
	 w_i = 24'b 111111111111111110000010;
	 next_valid = 1'b1;
	 end
	10'd727: begin 
	 w_r = 24'b 111111111111111100100000;
	 w_i = 24'b 111111111111111110000101;
	 next_valid = 1'b1;
	 end
	10'd728: begin 
	 w_r = 24'b 111111111111111100011110;
	 w_i = 24'b 111111111111111110000111;
	 next_valid = 1'b1;
	 end
	10'd729: begin 
	 w_r = 24'b 111111111111111100011101;
	 w_i = 24'b 111111111111111110001010;
	 next_valid = 1'b1;
	 end
	10'd730: begin 
	 w_r = 24'b 111111111111111100011011;
	 w_i = 24'b 111111111111111110001101;
	 next_valid = 1'b1;
	 end
	10'd731: begin 
	 w_r = 24'b 111111111111111100011010;
	 w_i = 24'b 111111111111111110010000;
	 next_valid = 1'b1;
	 end
	10'd732: begin 
	 w_r = 24'b 111111111111111100011001;
	 w_i = 24'b 111111111111111110010011;
	 next_valid = 1'b1;
	 end
	10'd733: begin 
	 w_r = 24'b 111111111111111100010111;
	 w_i = 24'b 111111111111111110010101;
	 next_valid = 1'b1;
	 end
	10'd734: begin 
	 w_r = 24'b 111111111111111100010110;
	 w_i = 24'b 111111111111111110011000;
	 next_valid = 1'b1;
	 end
	10'd735: begin 
	 w_r = 24'b 111111111111111100010101;
	 w_i = 24'b 111111111111111110011011;
	 next_valid = 1'b1;
	 end
	10'd736: begin 
	 w_r = 24'b 111111111111111100010011;
	 w_i = 24'b 111111111111111110011110;
	 next_valid = 1'b1;
	 end
	10'd737: begin 
	 w_r = 24'b 111111111111111100010010;
	 w_i = 24'b 111111111111111110100001;
	 next_valid = 1'b1;
	 end
	10'd738: begin 
	 w_r = 24'b 111111111111111100010001;
	 w_i = 24'b 111111111111111110100100;
	 next_valid = 1'b1;
	 end
	10'd739: begin 
	 w_r = 24'b 111111111111111100010000;
	 w_i = 24'b 111111111111111110100111;
	 next_valid = 1'b1;
	 end
	10'd740: begin 
	 w_r = 24'b 111111111111111100001111;
	 w_i = 24'b 111111111111111110101010;
	 next_valid = 1'b1;
	 end
	10'd741: begin 
	 w_r = 24'b 111111111111111100001110;
	 w_i = 24'b 111111111111111110101101;
	 next_valid = 1'b1;
	 end
	10'd742: begin 
	 w_r = 24'b 111111111111111100001101;
	 w_i = 24'b 111111111111111110110000;
	 next_valid = 1'b1;
	 end
	10'd743: begin 
	 w_r = 24'b 111111111111111100001100;
	 w_i = 24'b 111111111111111110110011;
	 next_valid = 1'b1;
	 end
	10'd744: begin 
	 w_r = 24'b 111111111111111100001011;
	 w_i = 24'b 111111111111111110110110;
	 next_valid = 1'b1;
	 end
	10'd745: begin 
	 w_r = 24'b 111111111111111100001010;
	 w_i = 24'b 111111111111111110111001;
	 next_valid = 1'b1;
	 end
	10'd746: begin 
	 w_r = 24'b 111111111111111100001001;
	 w_i = 24'b 111111111111111110111100;
	 next_valid = 1'b1;
	 end
	10'd747: begin 
	 w_r = 24'b 111111111111111100001000;
	 w_i = 24'b 111111111111111110111111;
	 next_valid = 1'b1;
	 end
	10'd748: begin 
	 w_r = 24'b 111111111111111100001000;
	 w_i = 24'b 111111111111111111000010;
	 next_valid = 1'b1;
	 end
	10'd749: begin 
	 w_r = 24'b 111111111111111100000111;
	 w_i = 24'b 111111111111111111000101;
	 next_valid = 1'b1;
	 end
	10'd750: begin 
	 w_r = 24'b 111111111111111100000110;
	 w_i = 24'b 111111111111111111001000;
	 next_valid = 1'b1;
	 end
	10'd751: begin 
	 w_r = 24'b 111111111111111100000110;
	 w_i = 24'b 111111111111111111001011;
	 next_valid = 1'b1;
	 end
	10'd752: begin 
	 w_r = 24'b 111111111111111100000101;
	 w_i = 24'b 111111111111111111001110;
	 next_valid = 1'b1;
	 end
	10'd753: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010001;
	 next_valid = 1'b1;
	 end
	10'd754: begin 
	 w_r = 24'b 111111111111111100000100;
	 w_i = 24'b 111111111111111111010100;
	 next_valid = 1'b1;
	 end
	10'd755: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111010111;
	 next_valid = 1'b1;
	 end
	10'd756: begin 
	 w_r = 24'b 111111111111111100000011;
	 w_i = 24'b 111111111111111111011010;
	 next_valid = 1'b1;
	 end
	10'd757: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111011110;
	 next_valid = 1'b1;
	 end
	10'd758: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111100001;
	 next_valid = 1'b1;
	 end
	10'd759: begin 
	 w_r = 24'b 111111111111111100000010;
	 w_i = 24'b 111111111111111111100100;
	 next_valid = 1'b1;
	 end
	10'd760: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111100111;
	 next_valid = 1'b1;
	 end
	10'd761: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101010;
	 next_valid = 1'b1;
	 end
	10'd762: begin 
	 w_r = 24'b 111111111111111100000001;
	 w_i = 24'b 111111111111111111101101;
	 next_valid = 1'b1;
	 end
	10'd763: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110000;
	 next_valid = 1'b1;
	 end
	10'd764: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110011;
	 next_valid = 1'b1;
	 end
	10'd765: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111110111;
	 next_valid = 1'b1;
	 end
	10'd766: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111010;
	 next_valid = 1'b1;
	 end
	10'd767: begin 
	 w_r = 24'b 111111111111111100000000;
	 w_i = 24'b 111111111111111111111101;
	 next_valid = 1'b0;
	 end
	default: begin 
	 w_r = 24'b 000000000000000100000000;
	 w_i = 24'b 000000000000000000000000;
	 next_valid = 1'b1;
	 end
	endcase
end
////////////////////////////////////////////
// State register
always@(posedge clk or negedge rst_n)begin
    if(~rst_n)begin
        count <= 0;
        valid <= 0;
    end
    else if(in_valid)
    begin
        count <= next_count;
        valid <= in_valid;
    end
    else if (valid)
    begin
        count <= next_count;
        valid <= next_valid;
    end
end
endmodule