module FFT512_tb;
	parameter 					FFT_size		= 512;
	parameter 					IN_width		= 12;
	parameter 					OUT_width		= 16;
	parameter 					latency_limit	= 1030;
	parameter 					cycle			= 10.0;
	integer 					j;
    reg signed	[IN_width-1:0]  int_r           [0:FFT_size-1];
    reg signed	[IN_width-1:0]  int_i           [0:FFT_size-1];
	reg 						clk, rst_n, in_valid;
	wire 						out_valid;
	reg signed  [IN_width-1:0] 	din_r, din_i;
	wire signed [OUT_width-1:0] dout_r, dout_i;
////////////////////////////////////////////
	always #(cycle/2.0) 
		clk = ~clk;
////////////////////////////////////////////
	FFT512 uut_FFT512(
		.clk(clk),
		.rst_n(rst_n),
		.in_valid(in_valid),
		.din_r(din_r),
		.din_i(din_i),
		.out_valid(out_valid),
		.dout_r(dout_r),
		.dout_i(dout_i)
	);
////////////////////////////////////////////	
	initial begin
		int_r[0] =  0;
		int_r[1] =  331;
		int_r[2] =  229;
		int_r[3] =  -21;
		int_r[4] =  92;
		int_r[5] =  437;
		int_r[6] =  450;
		int_r[7] =  90;
		int_r[8] =  -93;
		int_r[9] =  119;
		int_r[10] =  256;
		int_r[11] =  -40;
		int_r[12] =  -394;
		int_r[13] =  -324;
		int_r[14] =  -37;
		int_r[15] =  -75;
		int_r[16] =  -394;
		int_r[17] =  -436;
		int_r[18] =  -72;
		int_r[19] =  173;
		int_r[20] =  0;
		int_r[21] =  -174;
		int_r[22] =  71;
		int_r[23] =  435;
		int_r[24] =  393;
		int_r[25] =  74;
		int_r[26] =  36;
		int_r[27] =  323;
		int_r[28] =  393;
		int_r[29] =  39;
		int_r[30] =  -256;
		int_r[31] =  -120;
		int_r[32] =  92;
		int_r[33] =  -91;
		int_r[34] =  -451;
		int_r[35] =  -438;
		int_r[36] =  -93;
		int_r[37] =  20;
		int_r[38] =  -230;
		int_r[39] =  -332;
		int_r[40] =  -1;
		int_r[41] =  331;
		int_r[42] =  229;
		int_r[43] =  -21;
		int_r[44] =  92;
		int_r[45] =  437;
		int_r[46] =  450;
		int_r[47] =  90;
		int_r[48] =  -93;
		int_r[49] =  119;
		int_r[50] =  256;
		int_r[51] =  -40;
		int_r[52] =  -394;
		int_r[53] =  -324;
		int_r[54] =  -37;
		int_r[55] =  -75;
		int_r[56] =  -394;
		int_r[57] =  -436;
		int_r[58] =  -72;
		int_r[59] =  173;
		int_r[60] =  0;
		int_r[61] =  -174;
		int_r[62] =  71;
		int_r[63] =  435;
		int_r[64] =  393;
		int_r[65] =  74;
		int_r[66] =  36;
		int_r[67] =  323;
		int_r[68] =  393;
		int_r[69] =  39;
		int_r[70] =  -256;
		int_r[71] =  -120;
		int_r[72] =  92;
		int_r[73] =  -91;
		int_r[74] =  -451;
		int_r[75] =  -438;
		int_r[76] =  -93;
		int_r[77] =  20;
		int_r[78] =  -230;
		int_r[79] =  -332;
		int_r[80] =  -1;
		int_r[81] =  331;
		int_r[82] =  229;
		int_r[83] =  -21;
		int_r[84] =  92;
		int_r[85] =  437;
		int_r[86] =  450;
		int_r[87] =  90;
		int_r[88] =  -93;
		int_r[89] =  119;
		int_r[90] =  256;
		int_r[91] =  -40;
		int_r[92] =  -394;
		int_r[93] =  -324;
		int_r[94] =  -37;
		int_r[95] =  -75;
		int_r[96] =  -394;
		int_r[97] =  -436;
		int_r[98] =  -72;
		int_r[99] =  173;
		int_r[100] =  0;
		int_r[101] =  -174;
		int_r[102] =  71;
		int_r[103] =  435;
		int_r[104] =  393;
		int_r[105] =  74;
		int_r[106] =  36;
		int_r[107] =  323;
		int_r[108] =  393;
		int_r[109] =  39;
		int_r[110] =  -256;
		int_r[111] =  -120;
		int_r[112] =  92;
		int_r[113] =  -91;
		int_r[114] =  -451;
		int_r[115] =  -438;
		int_r[116] =  -93;
		int_r[117] =  20;
		int_r[118] =  -230;
		int_r[119] =  -332;
		int_r[120] =  -1;
		int_r[121] =  331;
		int_r[122] =  229;
		int_r[123] =  -21;
		int_r[124] =  92;
		int_r[125] =  437;
		int_r[126] =  450;
		int_r[127] =  90;
		int_r[128] =  -93;
		int_r[129] =  119;
		int_r[130] =  255;
		int_r[131] =  -40;
		int_r[132] =  -394;
		int_r[133] =  -324;
		int_r[134] =  -37;
		int_r[135] =  -75;
		int_r[136] =  -394;
		int_r[137] =  -436;
		int_r[138] =  -72;
		int_r[139] =  173;
		int_r[140] =  -1;
		int_r[141] =  -174;
		int_r[142] =  71;
		int_r[143] =  435;
		int_r[144] =  393;
		int_r[145] =  74;
		int_r[146] =  36;
		int_r[147] =  323;
		int_r[148] =  393;
		int_r[149] =  39;
		int_r[150] =  -256;
		int_r[151] =  -120;
		int_r[152] =  92;
		int_r[153] =  -91;
		int_r[154] =  -451;
		int_r[155] =  -438;
		int_r[156] =  -93;
		int_r[157] =  20;
		int_r[158] =  -230;
		int_r[159] =  -332;
		int_r[160] =  -1;
		int_r[161] =  331;
		int_r[162] =  229;
		int_r[163] =  -21;
		int_r[164] =  92;
		int_r[165] =  437;
		int_r[166] =  450;
		int_r[167] =  90;
		int_r[168] =  -93;
		int_r[169] =  119;
		int_r[170] =  255;
		int_r[171] =  -40;
		int_r[172] =  -394;
		int_r[173] =  -324;
		int_r[174] =  -37;
		int_r[175] =  -75;
		int_r[176] =  -394;
		int_r[177] =  -436;
		int_r[178] =  -72;
		int_r[179] =  173;
		int_r[180] =  0;
		int_r[181] =  -174;
		int_r[182] =  71;
		int_r[183] =  435;
		int_r[184] =  393;
		int_r[185] =  74;
		int_r[186] =  36;
		int_r[187] =  323;
		int_r[188] =  393;
		int_r[189] =  39;
		int_r[190] =  -256;
		int_r[191] =  -120;
		int_r[192] =  92;
		int_r[193] =  -91;
		int_r[194] =  -451;
		int_r[195] =  -438;
		int_r[196] =  -93;
		int_r[197] =  20;
		int_r[198] =  -230;
		int_r[199] =  -332;
		int_r[200] =  -1;
		int_r[201] =  331;
		int_r[202] =  229;
		int_r[203] =  -21;
		int_r[204] =  92;
		int_r[205] =  437;
		int_r[206] =  450;
		int_r[207] =  90;
		int_r[208] =  -93;
		int_r[209] =  119;
		int_r[210] =  255;
		int_r[211] =  -40;
		int_r[212] =  -394;
		int_r[213] =  -324;
		int_r[214] =  -37;
		int_r[215] =  -75;
		int_r[216] =  -394;
		int_r[217] =  -436;
		int_r[218] =  -72;
		int_r[219] =  173;
		int_r[220] =  -1;
		int_r[221] =  -174;
		int_r[222] =  71;
		int_r[223] =  435;
		int_r[224] =  393;
		int_r[225] =  74;
		int_r[226] =  36;
		int_r[227] =  323;
		int_r[228] =  393;
		int_r[229] =  39;
		int_r[230] =  -256;
		int_r[231] =  -120;
		int_r[232] =  92;
		int_r[233] =  -91;
		int_r[234] =  -451;
		int_r[235] =  -438;
		int_r[236] =  -93;
		int_r[237] =  20;
		int_r[238] =  -230;
		int_r[239] =  -332;
		int_r[240] =  -1;
		int_r[241] =  331;
		int_r[242] =  229;
		int_r[243] =  -21;
		int_r[244] =  92;
		int_r[245] =  437;
		int_r[246] =  450;
		int_r[247] =  90;
		int_r[248] =  -93;
		int_r[249] =  119;
		int_r[250] =  255;
		int_r[251] =  -40;
		int_r[252] =  -394;
		int_r[253] =  -324;
		int_r[254] =  -37;
		int_r[255] =  -75;
		int_r[256] =  -394;
		int_r[257] =  -436;
		int_r[258] =  -72;
		int_r[259] =  173;
		int_r[260] =  0;
		int_r[261] =  -174;
		int_r[262] =  71;
		int_r[263] =  435;
		int_r[264] =  393;
		int_r[265] =  74;
		int_r[266] =  36;
		int_r[267] =  323;
		int_r[268] =  393;
		int_r[269] =  39;
		int_r[270] =  -256;
		int_r[271] =  -120;
		int_r[272] =  92;
		int_r[273] =  -91;
		int_r[274] =  -451;
		int_r[275] =  -438;
		int_r[276] =  -93;
		int_r[277] =  20;
		int_r[278] =  -230;
		int_r[279] =  -332;
		int_r[280] =  0;
		int_r[281] =  331;
		int_r[282] =  229;
		int_r[283] =  -21;
		int_r[284] =  92;
		int_r[285] =  437;
		int_r[286] =  450;
		int_r[287] =  90;
		int_r[288] =  -93;
		int_r[289] =  119;
		int_r[290] =  256;
		int_r[291] =  -40;
		int_r[292] =  -394;
		int_r[293] =  -324;
		int_r[294] =  -37;
		int_r[295] =  -75;
		int_r[296] =  -394;
		int_r[297] =  -436;
		int_r[298] =  -72;
		int_r[299] =  173;
		int_r[300] =  0;
		int_r[301] =  -174;
		int_r[302] =  71;
		int_r[303] =  435;
		int_r[304] =  393;
		int_r[305] =  74;
		int_r[306] =  36;
		int_r[307] =  323;
		int_r[308] =  393;
		int_r[309] =  39;
		int_r[310] =  -256;
		int_r[311] =  -120;
		int_r[312] =  92;
		int_r[313] =  -91;
		int_r[314] =  -451;
		int_r[315] =  -438;
		int_r[316] =  -93;
		int_r[317] =  20;
		int_r[318] =  -230;
		int_r[319] =  -332;
		int_r[320] =  -1;
		int_r[321] =  331;
		int_r[322] =  229;
		int_r[323] =  -21;
		int_r[324] =  92;
		int_r[325] =  437;
		int_r[326] =  450;
		int_r[327] =  90;
		int_r[328] =  -93;
		int_r[329] =  119;
		int_r[330] =  256;
		int_r[331] =  -40;
		int_r[332] =  -394;
		int_r[333] =  -324;
		int_r[334] =  -37;
		int_r[335] =  -75;
		int_r[336] =  -394;
		int_r[337] =  -436;
		int_r[338] =  -72;
		int_r[339] =  173;
		int_r[340] =  0;
		int_r[341] =  -174;
		int_r[342] =  71;
		int_r[343] =  435;
		int_r[344] =  393;
		int_r[345] =  74;
		int_r[346] =  36;
		int_r[347] =  323;
		int_r[348] =  393;
		int_r[349] =  39;
		int_r[350] =  -256;
		int_r[351] =  -120;
		int_r[352] =  92;
		int_r[353] =  -91;
		int_r[354] =  -451;
		int_r[355] =  -438;
		int_r[356] =  -93;
		int_r[357] =  20;
		int_r[358] =  -230;
		int_r[359] =  -332;
		int_r[360] =  -1;
		int_r[361] =  331;
		int_r[362] =  229;
		int_r[363] =  -21;
		int_r[364] =  92;
		int_r[365] =  437;
		int_r[366] =  450;
		int_r[367] =  90;
		int_r[368] =  -93;
		int_r[369] =  119;
		int_r[370] =  256;
		int_r[371] =  -40;
		int_r[372] =  -394;
		int_r[373] =  -324;
		int_r[374] =  -37;
		int_r[375] =  -75;
		int_r[376] =  -394;
		int_r[377] =  -436;
		int_r[378] =  -72;
		int_r[379] =  173;
		int_r[380] =  0;
		int_r[381] =  -174;
		int_r[382] =  71;
		int_r[383] =  435;
		int_r[384] =  393;
		int_r[385] =  74;
		int_r[386] =  36;
		int_r[387] =  323;
		int_r[388] =  393;
		int_r[389] =  39;
		int_r[390] =  -256;
		int_r[391] =  -120;
		int_r[392] =  92;
		int_r[393] =  -91;
		int_r[394] =  -451;
		int_r[395] =  -438;
		int_r[396] =  -93;
		int_r[397] =  20;
		int_r[398] =  -230;
		int_r[399] =  -332;
		int_r[400] =  -1;
		int_r[401] =  331;
		int_r[402] =  229;
		int_r[403] =  -21;
		int_r[404] =  92;
		int_r[405] =  437;
		int_r[406] =  450;
		int_r[407] =  90;
		int_r[408] =  -93;
		int_r[409] =  119;
		int_r[410] =  256;
		int_r[411] =  -40;
		int_r[412] =  -394;
		int_r[413] =  -324;
		int_r[414] =  -37;
		int_r[415] =  -75;
		int_r[416] =  -394;
		int_r[417] =  -436;
		int_r[418] =  -72;
		int_r[419] =  173;
		int_r[420] =  -1;
		int_r[421] =  -174;
		int_r[422] =  71;
		int_r[423] =  435;
		int_r[424] =  393;
		int_r[425] =  74;
		int_r[426] =  36;
		int_r[427] =  323;
		int_r[428] =  393;
		int_r[429] =  39;
		int_r[430] =  -256;
		int_r[431] =  -120;
		int_r[432] =  92;
		int_r[433] =  -91;
		int_r[434] =  -451;
		int_r[435] =  -438;
		int_r[436] =  -93;
		int_r[437] =  20;
		int_r[438] =  -230;
		int_r[439] =  -332;
		int_r[440] =  0;
		int_r[441] =  331;
		int_r[442] =  229;
		int_r[443] =  -21;
		int_r[444] =  92;
		int_r[445] =  437;
		int_r[446] =  450;
		int_r[447] =  90;
		int_r[448] =  -93;
		int_r[449] =  119;
		int_r[450] =  256;
		int_r[451] =  -40;
		int_r[452] =  -394;
		int_r[453] =  -324;
		int_r[454] =  -37;
		int_r[455] =  -75;
		int_r[456] =  -394;
		int_r[457] =  -436;
		int_r[458] =  -72;
		int_r[459] =  173;
		int_r[460] =  0;
		int_r[461] =  -174;
		int_r[462] =  71;
		int_r[463] =  435;
		int_r[464] =  393;
		int_r[465] =  74;
		int_r[466] =  36;
		int_r[467] =  323;
		int_r[468] =  393;
		int_r[469] =  39;
		int_r[470] =  -257;
		int_r[471] =  -120;
		int_r[472] =  92;
		int_r[473] =  -91;
		int_r[474] =  -451;
		int_r[475] =  -438;
		int_r[476] =  -93;
		int_r[477] =  20;
		int_r[478] =  -230;
		int_r[479] =  -332;
		int_r[480] =  -1;
		int_r[481] =  331;
		int_r[482] =  229;
		int_r[483] =  -21;
		int_r[484] =  92;
		int_r[485] =  437;
		int_r[486] =  450;
		int_r[487] =  90;
		int_r[488] =  -93;
		int_r[489] =  119;
		int_r[490] =  256;
		int_r[491] =  -40;
		int_r[492] =  -394;
		int_r[493] =  -324;
		int_r[494] =  -37;
		int_r[495] =  -75;
		int_r[496] =  -394;
		int_r[497] =  -436;
		int_r[498] =  -72;
		int_r[499] =  173;
		int_r[500] =  0;
		int_r[501] =  -174;
		int_r[502] =  71;
		int_r[503] =  435;
		int_r[504] =  393;
		int_r[505] =  74;
		int_r[506] =  36;
		int_r[507] =  323;
		int_r[508] =  393;
		int_r[509] =  39;
		int_r[510] =  -256;
		int_r[511] =  -120;
	end
	initial begin
		int_i[0] =  0;
		int_i[1] =  0;
		int_i[2] =  0;
		int_i[3] =  0;
		int_i[4] =  0;
		int_i[5] =  0;
		int_i[6] =  0;
		int_i[7] =  0;
		int_i[8] =  0;
		int_i[9] =  0;
		int_i[10] =  0;
		int_i[11] =  0;
		int_i[12] =  0;
		int_i[13] =  0;
		int_i[14] =  0;
		int_i[15] =  0;
		int_i[16] =  0;
		int_i[17] =  0;
		int_i[18] =  0;
		int_i[19] =  0;
		int_i[20] =  0;
		int_i[21] =  0;
		int_i[22] =  0;
		int_i[23] =  0;
		int_i[24] =  0;
		int_i[25] =  0;
		int_i[26] =  0;
		int_i[27] =  0;
		int_i[28] =  0;
		int_i[29] =  0;
		int_i[30] =  0;
		int_i[31] =  0;
		int_i[32] =  0;
		int_i[33] =  0;
		int_i[34] =  0;
		int_i[35] =  0;
		int_i[36] =  0;
		int_i[37] =  0;
		int_i[38] =  0;
		int_i[39] =  0;
		int_i[40] =  0;
		int_i[41] =  0;
		int_i[42] =  0;
		int_i[43] =  0;
		int_i[44] =  0;
		int_i[45] =  0;
		int_i[46] =  0;
		int_i[47] =  0;
		int_i[48] =  0;
		int_i[49] =  0;
		int_i[50] =  0;
		int_i[51] =  0;
		int_i[52] =  0;
		int_i[53] =  0;
		int_i[54] =  0;
		int_i[55] =  0;
		int_i[56] =  0;
		int_i[57] =  0;
		int_i[58] =  0;
		int_i[59] =  0;
		int_i[60] =  0;
		int_i[61] =  0;
		int_i[62] =  0;
		int_i[63] =  0;
		int_i[64] =  0;
		int_i[65] =  0;
		int_i[66] =  0;
		int_i[67] =  0;
		int_i[68] =  0;
		int_i[69] =  0;
		int_i[70] =  0;
		int_i[71] =  0;
		int_i[72] =  0;
		int_i[73] =  0;
		int_i[74] =  0;
		int_i[75] =  0;
		int_i[76] =  0;
		int_i[77] =  0;
		int_i[78] =  0;
		int_i[79] =  0;
		int_i[80] =  0;
		int_i[81] =  0;
		int_i[82] =  0;
		int_i[83] =  0;
		int_i[84] =  0;
		int_i[85] =  0;
		int_i[86] =  0;
		int_i[87] =  0;
		int_i[88] =  0;
		int_i[89] =  0;
		int_i[90] =  0;
		int_i[91] =  0;
		int_i[92] =  0;
		int_i[93] =  0;
		int_i[94] =  0;
		int_i[95] =  0;
		int_i[96] =  0;
		int_i[97] =  0;
		int_i[98] =  0;
		int_i[99] =  0;
		int_i[100] =  0;
		int_i[101] =  0;
		int_i[102] =  0;
		int_i[103] =  0;
		int_i[104] =  0;
		int_i[105] =  0;
		int_i[106] =  0;
		int_i[107] =  0;
		int_i[108] =  0;
		int_i[109] =  0;
		int_i[110] =  0;
		int_i[111] =  0;
		int_i[112] =  0;
		int_i[113] =  0;
		int_i[114] =  0;
		int_i[115] =  0;
		int_i[116] =  0;
		int_i[117] =  0;
		int_i[118] =  0;
		int_i[119] =  0;
		int_i[120] =  0;
		int_i[121] =  0;
		int_i[122] =  0;
		int_i[123] =  0;
		int_i[124] =  0;
		int_i[125] =  0;
		int_i[126] =  0;
		int_i[127] =  0;
		int_i[128] =  0;
		int_i[129] =  0;
		int_i[130] =  0;
		int_i[131] =  0;
		int_i[132] =  0;
		int_i[133] =  0;
		int_i[134] =  0;
		int_i[135] =  0;
		int_i[136] =  0;
		int_i[137] =  0;
		int_i[138] =  0;
		int_i[139] =  0;
		int_i[140] =  0;
		int_i[141] =  0;
		int_i[142] =  0;
		int_i[143] =  0;
		int_i[144] =  0;
		int_i[145] =  0;
		int_i[146] =  0;
		int_i[147] =  0;
		int_i[148] =  0;
		int_i[149] =  0;
		int_i[150] =  0;
		int_i[151] =  0;
		int_i[152] =  0;
		int_i[153] =  0;
		int_i[154] =  0;
		int_i[155] =  0;
		int_i[156] =  0;
		int_i[157] =  0;
		int_i[158] =  0;
		int_i[159] =  0;
		int_i[160] =  0;
		int_i[161] =  0;
		int_i[162] =  0;
		int_i[163] =  0;
		int_i[164] =  0;
		int_i[165] =  0;
		int_i[166] =  0;
		int_i[167] =  0;
		int_i[168] =  0;
		int_i[169] =  0;
		int_i[170] =  0;
		int_i[171] =  0;
		int_i[172] =  0;
		int_i[173] =  0;
		int_i[174] =  0;
		int_i[175] =  0;
		int_i[176] =  0;
		int_i[177] =  0;
		int_i[178] =  0;
		int_i[179] =  0;
		int_i[180] =  0;
		int_i[181] =  0;
		int_i[182] =  0;
		int_i[183] =  0;
		int_i[184] =  0;
		int_i[185] =  0;
		int_i[186] =  0;
		int_i[187] =  0;
		int_i[188] =  0;
		int_i[189] =  0;
		int_i[190] =  0;
		int_i[191] =  0;
		int_i[192] =  0;
		int_i[193] =  0;
		int_i[194] =  0;
		int_i[195] =  0;
		int_i[196] =  0;
		int_i[197] =  0;
		int_i[198] =  0;
		int_i[199] =  0;
		int_i[200] =  0;
		int_i[201] =  0;
		int_i[202] =  0;
		int_i[203] =  0;
		int_i[204] =  0;
		int_i[205] =  0;
		int_i[206] =  0;
		int_i[207] =  0;
		int_i[208] =  0;
		int_i[209] =  0;
		int_i[210] =  0;
		int_i[211] =  0;
		int_i[212] =  0;
		int_i[213] =  0;
		int_i[214] =  0;
		int_i[215] =  0;
		int_i[216] =  0;
		int_i[217] =  0;
		int_i[218] =  0;
		int_i[219] =  0;
		int_i[220] =  0;
		int_i[221] =  0;
		int_i[222] =  0;
		int_i[223] =  0;
		int_i[224] =  0;
		int_i[225] =  0;
		int_i[226] =  0;
		int_i[227] =  0;
		int_i[228] =  0;
		int_i[229] =  0;
		int_i[230] =  0;
		int_i[231] =  0;
		int_i[232] =  0;
		int_i[233] =  0;
		int_i[234] =  0;
		int_i[235] =  0;
		int_i[236] =  0;
		int_i[237] =  0;
		int_i[238] =  0;
		int_i[239] =  0;
		int_i[240] =  0;
		int_i[241] =  0;
		int_i[242] =  0;
		int_i[243] =  0;
		int_i[244] =  0;
		int_i[245] =  0;
		int_i[246] =  0;
		int_i[247] =  0;
		int_i[248] =  0;
		int_i[249] =  0;
		int_i[250] =  0;
		int_i[251] =  0;
		int_i[252] =  0;
		int_i[253] =  0;
		int_i[254] =  0;
		int_i[255] =  0;
		int_i[256] =  0;
		int_i[257] =  0;
		int_i[258] =  0;
		int_i[259] =  0;
		int_i[260] =  0;
		int_i[261] =  0;
		int_i[262] =  0;
		int_i[263] =  0;
		int_i[264] =  0;
		int_i[265] =  0;
		int_i[266] =  0;
		int_i[267] =  0;
		int_i[268] =  0;
		int_i[269] =  0;
		int_i[270] =  0;
		int_i[271] =  0;
		int_i[272] =  0;
		int_i[273] =  0;
		int_i[274] =  0;
		int_i[275] =  0;
		int_i[276] =  0;
		int_i[277] =  0;
		int_i[278] =  0;
		int_i[279] =  0;
		int_i[280] =  0;
		int_i[281] =  0;
		int_i[282] =  0;
		int_i[283] =  0;
		int_i[284] =  0;
		int_i[285] =  0;
		int_i[286] =  0;
		int_i[287] =  0;
		int_i[288] =  0;
		int_i[289] =  0;
		int_i[290] =  0;
		int_i[291] =  0;
		int_i[292] =  0;
		int_i[293] =  0;
		int_i[294] =  0;
		int_i[295] =  0;
		int_i[296] =  0;
		int_i[297] =  0;
		int_i[298] =  0;
		int_i[299] =  0;
		int_i[300] =  0;
		int_i[301] =  0;
		int_i[302] =  0;
		int_i[303] =  0;
		int_i[304] =  0;
		int_i[305] =  0;
		int_i[306] =  0;
		int_i[307] =  0;
		int_i[308] =  0;
		int_i[309] =  0;
		int_i[310] =  0;
		int_i[311] =  0;
		int_i[312] =  0;
		int_i[313] =  0;
		int_i[314] =  0;
		int_i[315] =  0;
		int_i[316] =  0;
		int_i[317] =  0;
		int_i[318] =  0;
		int_i[319] =  0;
		int_i[320] =  0;
		int_i[321] =  0;
		int_i[322] =  0;
		int_i[323] =  0;
		int_i[324] =  0;
		int_i[325] =  0;
		int_i[326] =  0;
		int_i[327] =  0;
		int_i[328] =  0;
		int_i[329] =  0;
		int_i[330] =  0;
		int_i[331] =  0;
		int_i[332] =  0;
		int_i[333] =  0;
		int_i[334] =  0;
		int_i[335] =  0;
		int_i[336] =  0;
		int_i[337] =  0;
		int_i[338] =  0;
		int_i[339] =  0;
		int_i[340] =  0;
		int_i[341] =  0;
		int_i[342] =  0;
		int_i[343] =  0;
		int_i[344] =  0;
		int_i[345] =  0;
		int_i[346] =  0;
		int_i[347] =  0;
		int_i[348] =  0;
		int_i[349] =  0;
		int_i[350] =  0;
		int_i[351] =  0;
		int_i[352] =  0;
		int_i[353] =  0;
		int_i[354] =  0;
		int_i[355] =  0;
		int_i[356] =  0;
		int_i[357] =  0;
		int_i[358] =  0;
		int_i[359] =  0;
		int_i[360] =  0;
		int_i[361] =  0;
		int_i[362] =  0;
		int_i[363] =  0;
		int_i[364] =  0;
		int_i[365] =  0;
		int_i[366] =  0;
		int_i[367] =  0;
		int_i[368] =  0;
		int_i[369] =  0;
		int_i[370] =  0;
		int_i[371] =  0;
		int_i[372] =  0;
		int_i[373] =  0;
		int_i[374] =  0;
		int_i[375] =  0;
		int_i[376] =  0;
		int_i[377] =  0;
		int_i[378] =  0;
		int_i[379] =  0;
		int_i[380] =  0;
		int_i[381] =  0;
		int_i[382] =  0;
		int_i[383] =  0;
		int_i[384] =  0;
		int_i[385] =  0;
		int_i[386] =  0;
		int_i[387] =  0;
		int_i[388] =  0;
		int_i[389] =  0;
		int_i[390] =  0;
		int_i[391] =  0;
		int_i[392] =  0;
		int_i[393] =  0;
		int_i[394] =  0;
		int_i[395] =  0;
		int_i[396] =  0;
		int_i[397] =  0;
		int_i[398] =  0;
		int_i[399] =  0;
		int_i[400] =  0;
		int_i[401] =  0;
		int_i[402] =  0;
		int_i[403] =  0;
		int_i[404] =  0;
		int_i[405] =  0;
		int_i[406] =  0;
		int_i[407] =  0;
		int_i[408] =  0;
		int_i[409] =  0;
		int_i[410] =  0;
		int_i[411] =  0;
		int_i[412] =  0;
		int_i[413] =  0;
		int_i[414] =  0;
		int_i[415] =  0;
		int_i[416] =  0;
		int_i[417] =  0;
		int_i[418] =  0;
		int_i[419] =  0;
		int_i[420] =  0;
		int_i[421] =  0;
		int_i[422] =  0;
		int_i[423] =  0;
		int_i[424] =  0;
		int_i[425] =  0;
		int_i[426] =  0;
		int_i[427] =  0;
		int_i[428] =  0;
		int_i[429] =  0;
		int_i[430] =  0;
		int_i[431] =  0;
		int_i[432] =  0;
		int_i[433] =  0;
		int_i[434] =  0;
		int_i[435] =  0;
		int_i[436] =  0;
		int_i[437] =  0;
		int_i[438] =  0;
		int_i[439] =  0;
		int_i[440] =  0;
		int_i[441] =  0;
		int_i[442] =  0;
		int_i[443] =  0;
		int_i[444] =  0;
		int_i[445] =  0;
		int_i[446] =  0;
		int_i[447] =  0;
		int_i[448] =  0;
		int_i[449] =  0;
		int_i[450] =  0;
		int_i[451] =  0;
		int_i[452] =  0;
		int_i[453] =  0;
		int_i[454] =  0;
		int_i[455] =  0;
		int_i[456] =  0;
		int_i[457] =  0;
		int_i[458] =  0;
		int_i[459] =  0;
		int_i[460] =  0;
		int_i[461] =  0;
		int_i[462] =  0;
		int_i[463] =  0;
		int_i[464] =  0;
		int_i[465] =  0;
		int_i[466] =  0;
		int_i[467] =  0;
		int_i[468] =  0;
		int_i[469] =  0;
		int_i[470] =  0;
		int_i[471] =  0;
		int_i[472] =  0;
		int_i[473] =  0;
		int_i[474] =  0;
		int_i[475] =  0;
		int_i[476] =  0;
		int_i[477] =  0;
		int_i[478] =  0;
		int_i[479] =  0;
		int_i[480] =  0;
		int_i[481] =  0;
		int_i[482] =  0;
		int_i[483] =  0;
		int_i[484] =  0;
		int_i[485] =  0;
		int_i[486] =  0;
		int_i[487] =  0;
		int_i[488] =  0;
		int_i[489] =  0;
		int_i[490] =  0;
		int_i[491] =  0;
		int_i[492] =  0;
		int_i[493] =  0;
		int_i[494] =  0;
		int_i[495] =  0;
		int_i[496] =  0;
		int_i[497] =  0;
		int_i[498] =  0;
		int_i[499] =  0;
		int_i[500] =  0;
		int_i[501] =  0;
		int_i[502] =  0;
		int_i[503] =  0;
		int_i[504] =  0;
		int_i[505] =  0;
		int_i[506] =  0;
		int_i[507] =  0;
		int_i[508] =  0;
		int_i[509] =  0;
		int_i[510] =  0;
		int_i[511] =  0;
	end
////////////////////////////////////////////	
	initial begin
		clk = 0;
		rst_n = 1;
		in_valid = 0;
		@(negedge clk);
		@(negedge clk)	rst_n = 0;
		@(negedge clk)  rst_n = 1;
		@(negedge clk);
		////////////////////////
		for(j=0;j<FFT_size;j=j+1) begin
			@(negedge clk);
			in_valid 	= 1;
			din_r 		= int_r[j];
			din_i 		= int_i[j];
		end
		@(negedge clk) in_valid = 0;
		////////////////////////
		////////////////////////
		for(j=0;j<FFT_size;j=j+1) begin
			while(!out_valid) begin
				@(negedge clk); 
			end
		@(negedge clk);	
		end
		///////////////////////
		///////////////////////		
		$stop;
	end
endmodule
	

